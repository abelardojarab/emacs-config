Test netlist for Eldo & Spice mode

!---------------------------------------------------------------
!-- Project       : (X)emacs eldo & spice mode
!-- Circuit name  : test_netlist.cir
!---------------------------------------------------------------
!-- Designer(s)   : E. ROUAT <emmanuel.rouat@.wanadoo.fr>
!                 : G. VAN DER PLAS <geert_vanderplas@email.com>
!-- Library       : 
!-- Purpose       : Test for eldo and spice mode 
!-- Inputs        : 
!-- Outputs       : 
!-- Supplies      : 
!-- References    : 
!---------------------------------------------------------------
mn2 1 2 3 4 pmos l=10u w=1u 
mn1 1 2 3 4 nmos w='10u*wscale' l=1u $x=10u $l=1u $ test this doc $y=1u ?
Xaaa 1 2 3 4 5 6 FOO 
+ param: test=10f $ test for eldo
*+ couple=5 $ couple only for layla/mondriaan

! Note the difference between 'comments' and 'doc strings' :

* This is a 'commented out' line
! and this is a 'doc' string
$ and this is also a 'doc' string
* and a combination !of $both $ tested
* and a combination !of both tested
* and a 'combination' $of both tested

! You can comment out portions of text using #c/#e:

#c
.model MY_NMOS NMOS LEVEL=3 
+ VTO=1V UO=550 VMAX=2.0e5 
+ CGDO=0.4p CGBO=2.0e-10

.model MY_PMOS NMOS LEVEL=3 
+ VTO=-1V UO=230 VMAX=1.9e5 
+ CGDO=0.4p CGBO=2.0e-10
#e

! By using 'C-c C-c' you can 'toggle' between commented out portions
! of test - select the region that follows, type 'C-c C-c' (or use
! the '(Un)comment-region menu)' and see what happens:

! <select from here>

.param Rload=1MEG
.param Cload=1nF
*.param Rload=10MEG
* .param Cload=0.1nF

! <to here>

!--------------------------------------------------------------------
!	LIBRARIES 
!--------------------------------------------------------------------

! 'models.lib' should highlight when the moude pointer passes over it.
! This means you can load this file using the middle moude button (if
! the file exists)

.include models.lib
.lib key=typical models.lib


! Lets define some MOSFET models - these should appear in
! the 'Models' entry in the menu.

.model MY_NMOS NMOS LEVEL=3 
+ VTO=1V UO=550 VMAX=2.0e5 
+ CGDO=0.4p CGBO=2.0e-10

.model MY_PMOS NMOS LEVEL=3 
+ VTO=-1V UO=230 VMAX=1.9e5 
+ CGDO=0.4p CGBO=2.0e-10

! The following has a wrong syntax - note the fontification

.model 1WRONG_SYNTAX NMOS
+ LEVEL =2  


!--------------------------------------------------------------------
!	NETLIST 
!--------------------------------------------------------------------

! Lets define a subckt - a parametrised inverter

.SUBCKT FOO IN OUT VDD VSS param: W=5u L=0.5U
MP OUT IN VDD VDD MY_PMOS W={3*W} L={L}
MN OUT IN VSS! VSS! MY_NMOS W={W} L={L}
.ENDS FOO


! In the following instanciations, FOO should be highlighted

X1 1 2 3 4 FOO 
X2 1 2 3 4 FOO param: W=10u L=1u
X3 1 2 3 4 FOO ! comment

! Even in multi-line instanciations:
X4 1 2 3 4 
+ FOO param: W=10u L=1u
X5 1 2 
+ 3 4 FOO param: W=10u L=1u


! This one doesn't work - probably never will, in spice-mode it works
Xfail 1 2 3 4 
* commented line 
+ FOO param: W=10u L=1u


! FOO#1 is a valid name, but 1AOO1 isn't:

X6 1 2 3 4 FOO#1
X7 1 2 3 4 1AOO1


! net names
MN1 N1N28 N1N105 VSS VSS n W=1.056u L=0.185u 
+  AD=0.209P AS=0.122P PD=0.755U PS=0.280U 
+  NRD=0.297 NRS=0.160 
MM1I47N3 N1I471N25 N1N28 N1N37 VSS n W=0.440U L=0.180U 
+  AD=0.062P AS=0.209P PD=0.280U PS=0.755U 
+  NRD=0.315 NRS=0.370 
MM1I47N1 N1I471N6 N1N31 N1I471N25 VSS n W=0.440U L=0.180U 
+  AD=0.062P AS=0.062P PD=0.280U PS=0.280U 
+  NRD=0.315 NRS=0.315 
MM1I47N2 VSS RB N1I471N6 VSS n W=0.440U L=0.180U 
+  AD=0.405P AS=0.062P PD=2.280U PS=0.280U 
+  NRD=0.918 NRS=0.315 
MM1I120N VSS N1N37 N1N31 VSS n W=1.090U L=0.187U 
+  AD=0.377P AS=0.421P PD=0.960U PS=1.850U 
+  NRD=0.820 NRS=0.274 
MM1I139N3 N1I1391N26 N1N31 VSS VSS n W=1.199U L=0.187U 
+  AD=0.194P AS=0.377P PD=0.375U PS=0.960U 
+  NRD=0.142 NRS=0.764 
MM1I139N1 N1I1391N44 RB N1I1391N26 VSS n W=1.120U L=0.180U 
+  AD=0.157P AS=0.194P PD=0.280U PS=0.375U 
+  NRD=0.125 NRS=0.142 

!--------------------------------------------------------------------
!	SIMULATION OPTIONS 
!--------------------------------------------------------------------



.options STAT=1 SIMUDIV=10 !Status reports
.options noascii nomod engnot  
.options nowarn=240 nowarn=902 nowarn=123 
.options eps=1e-7 itol=1e-6 gmin=1e-16 analog 
.options nobound_phase paramfly inclib 
.width out=80 
.temp 27 

! Now some inputs and supplies

VDD VDD 0 DC 5V
VSS VSS 0 DC 0

VIN IN 0 Pulse(0 5 1us 0.1ns 0.1ns 10ns 20ns)

! Simulation cards - fontified in 'eldo-analysis-face' or 'spice-analysis-face'

.op
.tran 0.1us 10us 

! What will we look at? All 'output' cards are fontified 
! in font-lock-preprocessor-face:

.plot tran V(IN) V(OUT)
.plot tra V(OUT) ! Note wrong syntax
.probe I V

.extract tran AVERAGE(I(VDD)) 

.END

ytest opamp1 n1 n2

!--------------------------------------------------------------------
!	Changelog 
!--------------------------------------------------------------------

** Thu Apr 11 2002 Geert Van der Plas <geert_vanderplas@email.com>

**    - added spice mode remarks

* Thu Apr  5 2001 E. ROUAT (DAIS) <emmanuel.rouat@st.com>

    - File created


*** Local Variables:
*** mode:spice
*** End:
